-- Generated PORTMAP Stub File: Created by Capture FPGA Flow
-- Matches PCB component pinout with simulation model
-- Created Tuesday, March 08, 2022 16:27:20 ???? (?W?�??)

