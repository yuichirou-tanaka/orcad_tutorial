module TestMod();

endmodule